module FPU_normalization();

endmodule
