task automatic simulus_direct();
    
endtask //automatic

task automatic simulus_random(
    
);
    
endtask //automatic