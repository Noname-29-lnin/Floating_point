module CTR_center #()();

endmodule

