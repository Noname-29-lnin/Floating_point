module FPU_add_sub (
    input logic                 i_add_sub   , // i_add_sub = 0 (ADD) | = 1 (SUB)
    input logic [31:0]          i_32_a      ,
    input logic [31:0]          i_32_b      ,
    output logic [31:0]         o_32_s      ,
    output logic                o_ov_flag   ,
    output logic                o_un_flag    
);



endmodule
