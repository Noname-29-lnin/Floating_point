module FPU_rounding_hardware();

endmodule
