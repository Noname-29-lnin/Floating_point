//      // verilator_coverage annotation
        module MAN_ALU #(
            parameter NUM_OP    = 1 ,
            parameter SIZE_MAN  = 28
        )(
%000005     input logic [NUM_OP-1:0]    i_fpu_op        ,
%000001     input logic                 i_sign_max      ,
%000001     input logic                 i_sign_min      ,
%000000     input logic [SIZE_MAN-1:0]  i_man_max       ,
%000001     input logic [SIZE_MAN-1:0]  i_man_min       ,
%000001     output logic [SIZE_MAN-1:0] o_man_alu       ,
%000002     output logic                o_overflow       
        );
        
%000003 logic w_i_carry;
%000001 logic [SIZE_MAN-1:0] w_n_man_b;
%000003 logic [SIZE_MAN-1:0] w_i_man_b;
%000005 logic w_overflow;
        
        assign w_i_carry = i_fpu_op ? ~(i_sign_max ^ i_sign_min) : (i_sign_max ^ i_sign_min);
        assign w_n_man_b = ~(i_man_min);
        assign w_i_man_b = w_i_carry ? w_n_man_b : i_man_min;
        
        CLA_28bit ALU_SUB_UNIT (
            .i_carry        (w_i_carry),
            .i_data_a       (i_man_max),
            .i_data_b       (w_i_man_b),
            .o_sum          (o_man_alu),
            .o_carry        (w_overflow)
        );
        
        assign o_overflow = w_i_carry ? 1'b0 : w_overflow;
        
        endmodule
        
