module LOPD_unit #(
    parameter SIZE_NUM  = 24
)(
    input logic [SIZE_NUM-1:0]  i_data      ,
    output logic [SIZE_NUM-1:0] o_pos_one   ,
    output logic                o_zero_flag  
);



endmodule
