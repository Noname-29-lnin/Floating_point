module SUM_unit #(
    parameter SIZE_SUM  = 28
)();

endmodule