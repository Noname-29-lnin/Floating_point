module KSA_28bit(
    input logic         i_carry     ,
    input logic [27:0]  i_data_a    ,
    input logic [27:0]  i_data_b    ,
    output logic [27:0] o_sum       ,
    output logic        o_carry      
);


endmodule
