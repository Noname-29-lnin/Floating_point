module KSA_carry_graph #(
    parameter NUM_DEPTH     = 3 ,
    parameter SIZE_PADDED   = 8
)(
    input  logic [SIZE_PADDED-1:0]  i_p,
    input  logic [SIZE_PADDED-1:0]  i_g,
    output logic [SIZE_PADDED-1:0]  o_p,
    output logic [SIZE_PADDED-1:0]  o_g
);



endmodule
